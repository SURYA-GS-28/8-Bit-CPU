module instr_set (
    
);
    
endmodule